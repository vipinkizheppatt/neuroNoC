module PE(
	input a,
	input b,
	output c
);

always 
begin

end


endmodule